/***
Written by:  Nathan A. & Devin Nowowiejski
Date Written: 10-13-2025
Description: 3:1 Mux utilized throughout the SLP
cite:
	2:1 Multiplexer gotten from H&H, HDL Example 7.11 found on page 423
***/
module mux3 #(parameter WIDTH = 8)(
	input  logic [WIDTH-1:0] d0,
	input  logic [WIDTH-1:0] d1,
	input  logic [WIDTH-1:0] d2,
	input  logic [1:0]       s,
	output logic [WIDTH-1:0] y
);
	
	always_comb begin
		case (s)
			2'b00: y = d0;
			2'b01: y = d1;
			2'b10: y = d2;
			default: y = '0;
		endcase
	end
	
endmodule
