
/*
 * Written by: Brandon Kampsen & Luke Johnson
 * Date Written: 11-19-2025
 *
 * Description:
 *      This module is our conditional execution unit. It’s responsible for
 *      deciding whether an instruction is actually allowed to update anything
 *      (RegWrite, MemWrite, or PCSrc). We do this ARM-style: conditions are
 *      checked against the NZCV flags, and only if CondEx is true do we let
 *      the side-effects happen.
 *
 *      We also pipeline the flags in two halves (N/Z and C/V), just like the
 *      H&H example. That keeps the design simple and works well with our
 *      existing decode logic.
 */

module condunit
(

    // Basic clock + reset
    input  logic       CLK,           // main FPGA clock
    input  logic       reset,         // clears the flag registers

    // Condition + flag info
    input  logic [3:0] Cond,          // condition field from the instruction
    input  logic [3:0] ALUFlags,      // NZCV flags generated by ALU
    input  logic [1:0] FlagW,         // which halves of the flag register to update

    // Control signals that may or may not activate depending on CondEx
    input  logic       PCS,           // pipeline PCSrc control coming in
    input  logic       RegW,          // unconditioned register write enable
    input  logic       MemW,          // unconditioned memory write enable

    // Outputs after conditional gating
    output logic       PRSrc,         // conditioned PCSrc
    output logic       RegWrite,      // conditioned register write
    output logic       MemWrite       // conditioned data memory write
);

    logic [1:0] FlagWrite;   // determines which flag groups get updated
    logic [3:0] Flags;       // stored NZCV flags
    logic CondEx;            // whether the condition is satisfied


    // Flag register (split NZ / CV)
    flopenr #(2) flagreg_hi
	(
        .CLK(CLK),
        .reset(reset),
        .en(FlagWrite[1]),        // update N/Z if enabled
        .d(ALUFlags[3:2]),
        .q(Flags[3:2])
    );

    flopenr #(2) flagreg_lo
	(
        .CLK(CLK),
        .reset(reset),
        .en(FlagWrite[0]),        // update C/V if enabled
        .d(ALUFlags[1:0]),
        .q(Flags[1:0])
    );


    // Condition checking (ARM-style)
    condcheck cc
	(
        .Cond(Cond),
        .Flags(Flags),
        .CondEx(CondEx)
    );


    // ------------------------------
    // Conditional gating
    // ------------------------------
    assign FlagWrite = FlagW & {2{CondEx}};   // only write flags if condition passes
    assign RegWrite  = RegW  & CondEx;        // conditional register write
    assign MemWrite  = MemW  & CondEx;        // conditional memory write
    assign PRSrc     = PCS   & CondEx;        // conditional PC update

endmodule














/***
Written by:  Nathan A. & Devin Nowowiejski
Date Written: 11-3-2025
Description: Condiotional Unit for Pipeline Processor
cite: This Conditional Unit was found from H&H pg. 416, HDL Example 7.4
	Resettable Flip-Flop gotten from H&H, HDL Example 7.9 found on page 422
***/

// Add header 
/*
module condunit(
	input  logic       CLK,
	input  logic       reset,
	input  logic [3:0] Cond,
	input  logic [3:0] ALUFlags,
	input  logic [1:0] FlagW,
	input  logic       PCS,
	input  logic       RegW,
	input  logic       MemW,
	output logic       PRSrc,
	output logic       RegWrite,
	output logic       MemWrite
);
	logic [1:0] FlagWrite;
	logic [3:0] Flags;
	logic CondEx;

	// Split flag registers (N,Z) and (C,V)
	flopenr #(2) flagreg_hi(
		.CLK(CLK), .reset(reset), .en(FlagWrite[1]),
		.d(ALUFlags[3:2]), .q(Flags[3:2])
	);
	flopenr #(2) flagreg_lo(
		.CLK(CLK), .reset(reset), .en(FlagWrite[0]),
		.d(ALUFlags[1:0]), .q(Flags[1:0])
	);

	condcheck cc(
		.Cond(Cond),
		.Flags(Flags),
		.CondEx(CondEx)
	);

	assign FlagWrite = FlagW & {2{CondEx}};
	assign RegWrite  = RegW  & CondEx;
	assign MemWrite  = MemW  & CondEx;
	assign PRSrc     = PCS   & CondEx;
endmodule

*/


